module top;
bit signal_A;
bit signal_B; 
bit clk;


property chk;

endproperty


endmodule
