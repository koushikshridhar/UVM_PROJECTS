`include "uvm_pkg.sv"
import uvm_pkg::*;  //everything of uvm_pkg becomes part of my TB now

`include "mem_common.sv"
`include "memory.v"
`include "mem_tx.sv"
`include "mem_intf.sv"
`include "mem_reg_model.sv"
`include "mem_adaptor.sv"
`include "mem_sqr.sv"
`include "mem_drv.sv"
`include "seq_lib.sv"
`include "mem_agent.sv"
`include "mem_env.sv"
`include "test_lib.sv"
`include "top.sv"
